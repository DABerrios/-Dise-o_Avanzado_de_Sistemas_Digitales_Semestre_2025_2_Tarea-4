`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/06/2026 10:29:50 AM
// Design Name: 
// Module Name: coprocessor_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module coprocessor_top (
    input logic clk,      // 100 MHz System Clock
    input logic resetN,   // Reset 
    input logic rx,       // UART RX Pin
    output logic tx,      // UART TX Pin
    
    // --- Display Ports ---
    output logic [7:0] an,
    output logic [6:0] seg,
    output logic       dp
);

    // =========================================================================
    // SIGNALS
    // =========================================================================

    logic reset;
    assign reset = ~resetN; 

    clk_wiz_0 clkgen_i (
        .clk_in1      (clk),
        .reset        (~resetN),
        .clk_out1  (clk_out1),
        .locked       (wiz_locked)
    );
    
    logic [7:0] rx_data;
    logic       rx_ready;
    logic       tx_busy;
    logic       core_tx_start;
    logic [7:0] core_tx_data;

    logic       we_vec_1, we_vec_2;
    logic [9:0] mem_waddr;
    logic [9:0] mem_wdata;

    logic        ap_start;
    logic        ap_done, ap_ready, ap_idle;
    logic [47:0] hls_result;
    logic [1:0]  hls_opcode;

    logic [1023:0][9:0] q_A;
    logic [1023:0][9:0] q_B;
    
    logic [47:0] disp_data;
    logic [1:0]  disp_opcode;

    // =========================================================================
    // INSTANTIATIONS
    // =========================================================================

    // --- RX Control Logic
    rx_control ctrl_inst (
        .clk(clk_out1),
        .reset(reset), 
        .rx_data(rx_data), .rx_ready(rx_ready),
        .ap_done(ap_done), 
        .ap_start(ap_start), .hls_opcode(hls_opcode),
        .we_vec_1(we_vec_1), .we_vec_2(we_vec_2),
        .mem_waddr(mem_waddr), .mem_wdata(mem_wdata)
    );

    // --- memory
    wide_mem #(.TOTAL_ITEMS(1024)) mem_A (
        .clk(clk_out1),
        .wr_en(we_vec_1), .wr_addr(mem_waddr), .wr_data(mem_wdata), 
        .parallel_data(q_A) 
    );

    wide_mem #(.TOTAL_ITEMS(1024)) mem_B (
        .clk(clk_out1),
        .wr_en(we_vec_2), .wr_addr(mem_waddr), .wr_data(mem_wdata), 
        .parallel_data(q_B)
    );
    
    // --- core IP
    proc_core_0 hls_inst (
        .ap_clk(clk_out1),
        .ap_rst(reset), 
        .ap_start(ap_start),
        .ap_done(ap_done),
        .ap_idle(ap_idle),
        .ap_ready(ap_ready),
        .opcode(hls_opcode),
        .result(hls_result),
        
        .A_0(q_A[0]),
        .A_1(q_A[1]),
        .A_2(q_A[2]),
        .A_3(q_A[3]),
        .A_4(q_A[4]),
        .A_5(q_A[5]),
        .A_6(q_A[6]),
        .A_7(q_A[7]),
        .A_8(q_A[8]),
        .A_9(q_A[9]),
        .A_10(q_A[10]),
        .A_11(q_A[11]),
        .A_12(q_A[12]),
        .A_13(q_A[13]),
        .A_14(q_A[14]),
        .A_15(q_A[15]),
        .A_16(q_A[16]),
        .A_17(q_A[17]),
        .A_18(q_A[18]),
        .A_19(q_A[19]),
        .A_20(q_A[20]),
        .A_21(q_A[21]),
        .A_22(q_A[22]),
        .A_23(q_A[23]),
        .A_24(q_A[24]),
        .A_25(q_A[25]),
        .A_26(q_A[26]),
        .A_27(q_A[27]),
        .A_28(q_A[28]),
        .A_29(q_A[29]),
        .A_30(q_A[30]),
        .A_31(q_A[31]),
        .A_32(q_A[32]),
        .A_33(q_A[33]),
        .A_34(q_A[34]),
        .A_35(q_A[35]),
        .A_36(q_A[36]),
        .A_37(q_A[37]),
        .A_38(q_A[38]),
        .A_39(q_A[39]),
        .A_40(q_A[40]),
        .A_41(q_A[41]),
        .A_42(q_A[42]),
        .A_43(q_A[43]),
        .A_44(q_A[44]),
        .A_45(q_A[45]),
        .A_46(q_A[46]),
        .A_47(q_A[47]),
        .A_48(q_A[48]),
        .A_49(q_A[49]),
        .A_50(q_A[50]),
        .A_51(q_A[51]),
        .A_52(q_A[52]),
        .A_53(q_A[53]),
        .A_54(q_A[54]),
        .A_55(q_A[55]),
        .A_56(q_A[56]),
        .A_57(q_A[57]),
        .A_58(q_A[58]),
        .A_59(q_A[59]),
        .A_60(q_A[60]),
        .A_61(q_A[61]),
        .A_62(q_A[62]),
        .A_63(q_A[63]),
        .A_64(q_A[64]),
        .A_65(q_A[65]),
        .A_66(q_A[66]),
        .A_67(q_A[67]),
        .A_68(q_A[68]),
        .A_69(q_A[69]),
        .A_70(q_A[70]),
        .A_71(q_A[71]),
        .A_72(q_A[72]),
        .A_73(q_A[73]),
        .A_74(q_A[74]),
        .A_75(q_A[75]),
        .A_76(q_A[76]),
        .A_77(q_A[77]),
        .A_78(q_A[78]),
        .A_79(q_A[79]),
        .A_80(q_A[80]),
        .A_81(q_A[81]),
        .A_82(q_A[82]),
        .A_83(q_A[83]),
        .A_84(q_A[84]),
        .A_85(q_A[85]),
        .A_86(q_A[86]),
        .A_87(q_A[87]),
        .A_88(q_A[88]),
        .A_89(q_A[89]),
        .A_90(q_A[90]),
        .A_91(q_A[91]),
        .A_92(q_A[92]),
        .A_93(q_A[93]),
        .A_94(q_A[94]),
        .A_95(q_A[95]),
        .A_96(q_A[96]),
        .A_97(q_A[97]),
        .A_98(q_A[98]),
        .A_99(q_A[99]),
        .A_100(q_A[100]),
        .A_101(q_A[101]),
        .A_102(q_A[102]),
        .A_103(q_A[103]),
        .A_104(q_A[104]),
        .A_105(q_A[105]),
        .A_106(q_A[106]),
        .A_107(q_A[107]),
        .A_108(q_A[108]),
        .A_109(q_A[109]),
        .A_110(q_A[110]),
        .A_111(q_A[111]),
        .A_112(q_A[112]),
        .A_113(q_A[113]),
        .A_114(q_A[114]),
        .A_115(q_A[115]),
        .A_116(q_A[116]),
        .A_117(q_A[117]),
        .A_118(q_A[118]),
        .A_119(q_A[119]),
        .A_120(q_A[120]),
        .A_121(q_A[121]),
        .A_122(q_A[122]),
        .A_123(q_A[123]),
        .A_124(q_A[124]),
        .A_125(q_A[125]),
        .A_126(q_A[126]),
        .A_127(q_A[127]),
        .A_128(q_A[128]),
        .A_129(q_A[129]),
        .A_130(q_A[130]),
        .A_131(q_A[131]),
        .A_132(q_A[132]),
        .A_133(q_A[133]),
        .A_134(q_A[134]),
        .A_135(q_A[135]),
        .A_136(q_A[136]),
        .A_137(q_A[137]),
        .A_138(q_A[138]),
        .A_139(q_A[139]),
        .A_140(q_A[140]),
        .A_141(q_A[141]),
        .A_142(q_A[142]),
        .A_143(q_A[143]),
        .A_144(q_A[144]),
        .A_145(q_A[145]),
        .A_146(q_A[146]),
        .A_147(q_A[147]),
        .A_148(q_A[148]),
        .A_149(q_A[149]),
        .A_150(q_A[150]),
        .A_151(q_A[151]),
        .A_152(q_A[152]),
        .A_153(q_A[153]),
        .A_154(q_A[154]),
        .A_155(q_A[155]),
        .A_156(q_A[156]),
        .A_157(q_A[157]),
        .A_158(q_A[158]),
        .A_159(q_A[159]),
        .A_160(q_A[160]),
        .A_161(q_A[161]),
        .A_162(q_A[162]),
        .A_163(q_A[163]),
        .A_164(q_A[164]),
        .A_165(q_A[165]),
        .A_166(q_A[166]),
        .A_167(q_A[167]),
        .A_168(q_A[168]),
        .A_169(q_A[169]),
        .A_170(q_A[170]),
        .A_171(q_A[171]),
        .A_172(q_A[172]),
        .A_173(q_A[173]),
        .A_174(q_A[174]),
        .A_175(q_A[175]),
        .A_176(q_A[176]),
        .A_177(q_A[177]),
        .A_178(q_A[178]),
        .A_179(q_A[179]),
        .A_180(q_A[180]),
        .A_181(q_A[181]),
        .A_182(q_A[182]),
        .A_183(q_A[183]),
        .A_184(q_A[184]),
        .A_185(q_A[185]),
        .A_186(q_A[186]),
        .A_187(q_A[187]),
        .A_188(q_A[188]),
        .A_189(q_A[189]),
        .A_190(q_A[190]),
        .A_191(q_A[191]),
        .A_192(q_A[192]),
        .A_193(q_A[193]),
        .A_194(q_A[194]),
        .A_195(q_A[195]),
        .A_196(q_A[196]),
        .A_197(q_A[197]),
        .A_198(q_A[198]),
        .A_199(q_A[199]),
        .A_200(q_A[200]),
        .A_201(q_A[201]),
        .A_202(q_A[202]),
        .A_203(q_A[203]),
        .A_204(q_A[204]),
        .A_205(q_A[205]),
        .A_206(q_A[206]),
        .A_207(q_A[207]),
        .A_208(q_A[208]),
        .A_209(q_A[209]),
        .A_210(q_A[210]),
        .A_211(q_A[211]),
        .A_212(q_A[212]),
        .A_213(q_A[213]),
        .A_214(q_A[214]),
        .A_215(q_A[215]),
        .A_216(q_A[216]),
        .A_217(q_A[217]),
        .A_218(q_A[218]),
        .A_219(q_A[219]),
        .A_220(q_A[220]),
        .A_221(q_A[221]),
        .A_222(q_A[222]),
        .A_223(q_A[223]),
        .A_224(q_A[224]),
        .A_225(q_A[225]),
        .A_226(q_A[226]),
        .A_227(q_A[227]),
        .A_228(q_A[228]),
        .A_229(q_A[229]),
        .A_230(q_A[230]),
        .A_231(q_A[231]),
        .A_232(q_A[232]),
        .A_233(q_A[233]),
        .A_234(q_A[234]),
        .A_235(q_A[235]),
        .A_236(q_A[236]),
        .A_237(q_A[237]),
        .A_238(q_A[238]),
        .A_239(q_A[239]),
        .A_240(q_A[240]),
        .A_241(q_A[241]),
        .A_242(q_A[242]),
        .A_243(q_A[243]),
        .A_244(q_A[244]),
        .A_245(q_A[245]),
        .A_246(q_A[246]),
        .A_247(q_A[247]),
        .A_248(q_A[248]),
        .A_249(q_A[249]),
        .A_250(q_A[250]),
        .A_251(q_A[251]),
        .A_252(q_A[252]),
        .A_253(q_A[253]),
        .A_254(q_A[254]),
        .A_255(q_A[255]),
        .A_256(q_A[256]),
        .A_257(q_A[257]),
        .A_258(q_A[258]),
        .A_259(q_A[259]),
        .A_260(q_A[260]),
        .A_261(q_A[261]),
        .A_262(q_A[262]),
        .A_263(q_A[263]),
        .A_264(q_A[264]),
        .A_265(q_A[265]),
        .A_266(q_A[266]),
        .A_267(q_A[267]),
        .A_268(q_A[268]),
        .A_269(q_A[269]),
        .A_270(q_A[270]),
        .A_271(q_A[271]),
        .A_272(q_A[272]),
        .A_273(q_A[273]),
        .A_274(q_A[274]),
        .A_275(q_A[275]),
        .A_276(q_A[276]),
        .A_277(q_A[277]),
        .A_278(q_A[278]),
        .A_279(q_A[279]),
        .A_280(q_A[280]),
        .A_281(q_A[281]),
        .A_282(q_A[282]),
        .A_283(q_A[283]),
        .A_284(q_A[284]),
        .A_285(q_A[285]),
        .A_286(q_A[286]),
        .A_287(q_A[287]),
        .A_288(q_A[288]),
        .A_289(q_A[289]),
        .A_290(q_A[290]),
        .A_291(q_A[291]),
        .A_292(q_A[292]),
        .A_293(q_A[293]),
        .A_294(q_A[294]),
        .A_295(q_A[295]),
        .A_296(q_A[296]),
        .A_297(q_A[297]),
        .A_298(q_A[298]),
        .A_299(q_A[299]),
        .A_300(q_A[300]),
        .A_301(q_A[301]),
        .A_302(q_A[302]),
        .A_303(q_A[303]),
        .A_304(q_A[304]),
        .A_305(q_A[305]),
        .A_306(q_A[306]),
        .A_307(q_A[307]),
        .A_308(q_A[308]),
        .A_309(q_A[309]),
        .A_310(q_A[310]),
        .A_311(q_A[311]),
        .A_312(q_A[312]),
        .A_313(q_A[313]),
        .A_314(q_A[314]),
        .A_315(q_A[315]),
        .A_316(q_A[316]),
        .A_317(q_A[317]),
        .A_318(q_A[318]),
        .A_319(q_A[319]),
        .A_320(q_A[320]),
        .A_321(q_A[321]),
        .A_322(q_A[322]),
        .A_323(q_A[323]),
        .A_324(q_A[324]),
        .A_325(q_A[325]),
        .A_326(q_A[326]),
        .A_327(q_A[327]),
        .A_328(q_A[328]),
        .A_329(q_A[329]),
        .A_330(q_A[330]),
        .A_331(q_A[331]),
        .A_332(q_A[332]),
        .A_333(q_A[333]),
        .A_334(q_A[334]),
        .A_335(q_A[335]),
        .A_336(q_A[336]),
        .A_337(q_A[337]),
        .A_338(q_A[338]),
        .A_339(q_A[339]),
        .A_340(q_A[340]),
        .A_341(q_A[341]),
        .A_342(q_A[342]),
        .A_343(q_A[343]),
        .A_344(q_A[344]),
        .A_345(q_A[345]),
        .A_346(q_A[346]),
        .A_347(q_A[347]),
        .A_348(q_A[348]),
        .A_349(q_A[349]),
        .A_350(q_A[350]),
        .A_351(q_A[351]),
        .A_352(q_A[352]),
        .A_353(q_A[353]),
        .A_354(q_A[354]),
        .A_355(q_A[355]),
        .A_356(q_A[356]),
        .A_357(q_A[357]),
        .A_358(q_A[358]),
        .A_359(q_A[359]),
        .A_360(q_A[360]),
        .A_361(q_A[361]),
        .A_362(q_A[362]),
        .A_363(q_A[363]),
        .A_364(q_A[364]),
        .A_365(q_A[365]),
        .A_366(q_A[366]),
        .A_367(q_A[367]),
        .A_368(q_A[368]),
        .A_369(q_A[369]),
        .A_370(q_A[370]),
        .A_371(q_A[371]),
        .A_372(q_A[372]),
        .A_373(q_A[373]),
        .A_374(q_A[374]),
        .A_375(q_A[375]),
        .A_376(q_A[376]),
        .A_377(q_A[377]),
        .A_378(q_A[378]),
        .A_379(q_A[379]),
        .A_380(q_A[380]),
        .A_381(q_A[381]),
        .A_382(q_A[382]),
        .A_383(q_A[383]),
        .A_384(q_A[384]),
        .A_385(q_A[385]),
        .A_386(q_A[386]),
        .A_387(q_A[387]),
        .A_388(q_A[388]),
        .A_389(q_A[389]),
        .A_390(q_A[390]),
        .A_391(q_A[391]),
        .A_392(q_A[392]),
        .A_393(q_A[393]),
        .A_394(q_A[394]),
        .A_395(q_A[395]),
        .A_396(q_A[396]),
        .A_397(q_A[397]),
        .A_398(q_A[398]),
        .A_399(q_A[399]),
        .A_400(q_A[400]),
        .A_401(q_A[401]),
        .A_402(q_A[402]),
        .A_403(q_A[403]),
        .A_404(q_A[404]),
        .A_405(q_A[405]),
        .A_406(q_A[406]),
        .A_407(q_A[407]),
        .A_408(q_A[408]),
        .A_409(q_A[409]),
        .A_410(q_A[410]),
        .A_411(q_A[411]),
        .A_412(q_A[412]),
        .A_413(q_A[413]),
        .A_414(q_A[414]),
        .A_415(q_A[415]),
        .A_416(q_A[416]),
        .A_417(q_A[417]),
        .A_418(q_A[418]),
        .A_419(q_A[419]),
        .A_420(q_A[420]),
        .A_421(q_A[421]),
        .A_422(q_A[422]),
        .A_423(q_A[423]),
        .A_424(q_A[424]),
        .A_425(q_A[425]),
        .A_426(q_A[426]),
        .A_427(q_A[427]),
        .A_428(q_A[428]),
        .A_429(q_A[429]),
        .A_430(q_A[430]),
        .A_431(q_A[431]),
        .A_432(q_A[432]),
        .A_433(q_A[433]),
        .A_434(q_A[434]),
        .A_435(q_A[435]),
        .A_436(q_A[436]),
        .A_437(q_A[437]),
        .A_438(q_A[438]),
        .A_439(q_A[439]),
        .A_440(q_A[440]),
        .A_441(q_A[441]),
        .A_442(q_A[442]),
        .A_443(q_A[443]),
        .A_444(q_A[444]),
        .A_445(q_A[445]),
        .A_446(q_A[446]),
        .A_447(q_A[447]),
        .A_448(q_A[448]),
        .A_449(q_A[449]),
        .A_450(q_A[450]),
        .A_451(q_A[451]),
        .A_452(q_A[452]),
        .A_453(q_A[453]),
        .A_454(q_A[454]),
        .A_455(q_A[455]),
        .A_456(q_A[456]),
        .A_457(q_A[457]),
        .A_458(q_A[458]),
        .A_459(q_A[459]),
        .A_460(q_A[460]),
        .A_461(q_A[461]),
        .A_462(q_A[462]),
        .A_463(q_A[463]),
        .A_464(q_A[464]),
        .A_465(q_A[465]),
        .A_466(q_A[466]),
        .A_467(q_A[467]),
        .A_468(q_A[468]),
        .A_469(q_A[469]),
        .A_470(q_A[470]),
        .A_471(q_A[471]),
        .A_472(q_A[472]),
        .A_473(q_A[473]),
        .A_474(q_A[474]),
        .A_475(q_A[475]),
        .A_476(q_A[476]),
        .A_477(q_A[477]),
        .A_478(q_A[478]),
        .A_479(q_A[479]),
        .A_480(q_A[480]),
        .A_481(q_A[481]),
        .A_482(q_A[482]),
        .A_483(q_A[483]),
        .A_484(q_A[484]),
        .A_485(q_A[485]),
        .A_486(q_A[486]),
        .A_487(q_A[487]),
        .A_488(q_A[488]),
        .A_489(q_A[489]),
        .A_490(q_A[490]),
        .A_491(q_A[491]),
        .A_492(q_A[492]),
        .A_493(q_A[493]),
        .A_494(q_A[494]),
        .A_495(q_A[495]),
        .A_496(q_A[496]),
        .A_497(q_A[497]),
        .A_498(q_A[498]),
        .A_499(q_A[499]),
        .A_500(q_A[500]),
        .A_501(q_A[501]),
        .A_502(q_A[502]),
        .A_503(q_A[503]),
        .A_504(q_A[504]),
        .A_505(q_A[505]),
        .A_506(q_A[506]),
        .A_507(q_A[507]),
        .A_508(q_A[508]),
        .A_509(q_A[509]),
        .A_510(q_A[510]),
        .A_511(q_A[511]),
        .A_512(q_A[512]),
        .A_513(q_A[513]),
        .A_514(q_A[514]),
        .A_515(q_A[515]),
        .A_516(q_A[516]),
        .A_517(q_A[517]),
        .A_518(q_A[518]),
        .A_519(q_A[519]),
        .A_520(q_A[520]),
        .A_521(q_A[521]),
        .A_522(q_A[522]),
        .A_523(q_A[523]),
        .A_524(q_A[524]),
        .A_525(q_A[525]),
        .A_526(q_A[526]),
        .A_527(q_A[527]),
        .A_528(q_A[528]),
        .A_529(q_A[529]),
        .A_530(q_A[530]),
        .A_531(q_A[531]),
        .A_532(q_A[532]),
        .A_533(q_A[533]),
        .A_534(q_A[534]),
        .A_535(q_A[535]),
        .A_536(q_A[536]),
        .A_537(q_A[537]),
        .A_538(q_A[538]),
        .A_539(q_A[539]),
        .A_540(q_A[540]),
        .A_541(q_A[541]),
        .A_542(q_A[542]),
        .A_543(q_A[543]),
        .A_544(q_A[544]),
        .A_545(q_A[545]),
        .A_546(q_A[546]),
        .A_547(q_A[547]),
        .A_548(q_A[548]),
        .A_549(q_A[549]),
        .A_550(q_A[550]),
        .A_551(q_A[551]),
        .A_552(q_A[552]),
        .A_553(q_A[553]),
        .A_554(q_A[554]),
        .A_555(q_A[555]),
        .A_556(q_A[556]),
        .A_557(q_A[557]),
        .A_558(q_A[558]),
        .A_559(q_A[559]),
        .A_560(q_A[560]),
        .A_561(q_A[561]),
        .A_562(q_A[562]),
        .A_563(q_A[563]),
        .A_564(q_A[564]),
        .A_565(q_A[565]),
        .A_566(q_A[566]),
        .A_567(q_A[567]),
        .A_568(q_A[568]),
        .A_569(q_A[569]),
        .A_570(q_A[570]),
        .A_571(q_A[571]),
        .A_572(q_A[572]),
        .A_573(q_A[573]),
        .A_574(q_A[574]),
        .A_575(q_A[575]),
        .A_576(q_A[576]),
        .A_577(q_A[577]),
        .A_578(q_A[578]),
        .A_579(q_A[579]),
        .A_580(q_A[580]),
        .A_581(q_A[581]),
        .A_582(q_A[582]),
        .A_583(q_A[583]),
        .A_584(q_A[584]),
        .A_585(q_A[585]),
        .A_586(q_A[586]),
        .A_587(q_A[587]),
        .A_588(q_A[588]),
        .A_589(q_A[589]),
        .A_590(q_A[590]),
        .A_591(q_A[591]),
        .A_592(q_A[592]),
        .A_593(q_A[593]),
        .A_594(q_A[594]),
        .A_595(q_A[595]),
        .A_596(q_A[596]),
        .A_597(q_A[597]),
        .A_598(q_A[598]),
        .A_599(q_A[599]),
        .A_600(q_A[600]),
        .A_601(q_A[601]),
        .A_602(q_A[602]),
        .A_603(q_A[603]),
        .A_604(q_A[604]),
        .A_605(q_A[605]),
        .A_606(q_A[606]),
        .A_607(q_A[607]),
        .A_608(q_A[608]),
        .A_609(q_A[609]),
        .A_610(q_A[610]),
        .A_611(q_A[611]),
        .A_612(q_A[612]),
        .A_613(q_A[613]),
        .A_614(q_A[614]),
        .A_615(q_A[615]),
        .A_616(q_A[616]),
        .A_617(q_A[617]),
        .A_618(q_A[618]),
        .A_619(q_A[619]),
        .A_620(q_A[620]),
        .A_621(q_A[621]),
        .A_622(q_A[622]),
        .A_623(q_A[623]),
        .A_624(q_A[624]),
        .A_625(q_A[625]),
        .A_626(q_A[626]),
        .A_627(q_A[627]),
        .A_628(q_A[628]),
        .A_629(q_A[629]),
        .A_630(q_A[630]),
        .A_631(q_A[631]),
        .A_632(q_A[632]),
        .A_633(q_A[633]),
        .A_634(q_A[634]),
        .A_635(q_A[635]),
        .A_636(q_A[636]),
        .A_637(q_A[637]),
        .A_638(q_A[638]),
        .A_639(q_A[639]),
        .A_640(q_A[640]),
        .A_641(q_A[641]),
        .A_642(q_A[642]),
        .A_643(q_A[643]),
        .A_644(q_A[644]),
        .A_645(q_A[645]),
        .A_646(q_A[646]),
        .A_647(q_A[647]),
        .A_648(q_A[648]),
        .A_649(q_A[649]),
        .A_650(q_A[650]),
        .A_651(q_A[651]),
        .A_652(q_A[652]),
        .A_653(q_A[653]),
        .A_654(q_A[654]),
        .A_655(q_A[655]),
        .A_656(q_A[656]),
        .A_657(q_A[657]),
        .A_658(q_A[658]),
        .A_659(q_A[659]),
        .A_660(q_A[660]),
        .A_661(q_A[661]),
        .A_662(q_A[662]),
        .A_663(q_A[663]),
        .A_664(q_A[664]),
        .A_665(q_A[665]),
        .A_666(q_A[666]),
        .A_667(q_A[667]),
        .A_668(q_A[668]),
        .A_669(q_A[669]),
        .A_670(q_A[670]),
        .A_671(q_A[671]),
        .A_672(q_A[672]),
        .A_673(q_A[673]),
        .A_674(q_A[674]),
        .A_675(q_A[675]),
        .A_676(q_A[676]),
        .A_677(q_A[677]),
        .A_678(q_A[678]),
        .A_679(q_A[679]),
        .A_680(q_A[680]),
        .A_681(q_A[681]),
        .A_682(q_A[682]),
        .A_683(q_A[683]),
        .A_684(q_A[684]),
        .A_685(q_A[685]),
        .A_686(q_A[686]),
        .A_687(q_A[687]),
        .A_688(q_A[688]),
        .A_689(q_A[689]),
        .A_690(q_A[690]),
        .A_691(q_A[691]),
        .A_692(q_A[692]),
        .A_693(q_A[693]),
        .A_694(q_A[694]),
        .A_695(q_A[695]),
        .A_696(q_A[696]),
        .A_697(q_A[697]),
        .A_698(q_A[698]),
        .A_699(q_A[699]),
        .A_700(q_A[700]),
        .A_701(q_A[701]),
        .A_702(q_A[702]),
        .A_703(q_A[703]),
        .A_704(q_A[704]),
        .A_705(q_A[705]),
        .A_706(q_A[706]),
        .A_707(q_A[707]),
        .A_708(q_A[708]),
        .A_709(q_A[709]),
        .A_710(q_A[710]),
        .A_711(q_A[711]),
        .A_712(q_A[712]),
        .A_713(q_A[713]),
        .A_714(q_A[714]),
        .A_715(q_A[715]),
        .A_716(q_A[716]),
        .A_717(q_A[717]),
        .A_718(q_A[718]),
        .A_719(q_A[719]),
        .A_720(q_A[720]),
        .A_721(q_A[721]),
        .A_722(q_A[722]),
        .A_723(q_A[723]),
        .A_724(q_A[724]),
        .A_725(q_A[725]),
        .A_726(q_A[726]),
        .A_727(q_A[727]),
        .A_728(q_A[728]),
        .A_729(q_A[729]),
        .A_730(q_A[730]),
        .A_731(q_A[731]),
        .A_732(q_A[732]),
        .A_733(q_A[733]),
        .A_734(q_A[734]),
        .A_735(q_A[735]),
        .A_736(q_A[736]),
        .A_737(q_A[737]),
        .A_738(q_A[738]),
        .A_739(q_A[739]),
        .A_740(q_A[740]),
        .A_741(q_A[741]),
        .A_742(q_A[742]),
        .A_743(q_A[743]),
        .A_744(q_A[744]),
        .A_745(q_A[745]),
        .A_746(q_A[746]),
        .A_747(q_A[747]),
        .A_748(q_A[748]),
        .A_749(q_A[749]),
        .A_750(q_A[750]),
        .A_751(q_A[751]),
        .A_752(q_A[752]),
        .A_753(q_A[753]),
        .A_754(q_A[754]),
        .A_755(q_A[755]),
        .A_756(q_A[756]),
        .A_757(q_A[757]),
        .A_758(q_A[758]),
        .A_759(q_A[759]),
        .A_760(q_A[760]),
        .A_761(q_A[761]),
        .A_762(q_A[762]),
        .A_763(q_A[763]),
        .A_764(q_A[764]),
        .A_765(q_A[765]),
        .A_766(q_A[766]),
        .A_767(q_A[767]),
        .A_768(q_A[768]),
        .A_769(q_A[769]),
        .A_770(q_A[770]),
        .A_771(q_A[771]),
        .A_772(q_A[772]),
        .A_773(q_A[773]),
        .A_774(q_A[774]),
        .A_775(q_A[775]),
        .A_776(q_A[776]),
        .A_777(q_A[777]),
        .A_778(q_A[778]),
        .A_779(q_A[779]),
        .A_780(q_A[780]),
        .A_781(q_A[781]),
        .A_782(q_A[782]),
        .A_783(q_A[783]),
        .A_784(q_A[784]),
        .A_785(q_A[785]),
        .A_786(q_A[786]),
        .A_787(q_A[787]),
        .A_788(q_A[788]),
        .A_789(q_A[789]),
        .A_790(q_A[790]),
        .A_791(q_A[791]),
        .A_792(q_A[792]),
        .A_793(q_A[793]),
        .A_794(q_A[794]),
        .A_795(q_A[795]),
        .A_796(q_A[796]),
        .A_797(q_A[797]),
        .A_798(q_A[798]),
        .A_799(q_A[799]),
        .A_800(q_A[800]),
        .A_801(q_A[801]),
        .A_802(q_A[802]),
        .A_803(q_A[803]),
        .A_804(q_A[804]),
        .A_805(q_A[805]),
        .A_806(q_A[806]),
        .A_807(q_A[807]),
        .A_808(q_A[808]),
        .A_809(q_A[809]),
        .A_810(q_A[810]),
        .A_811(q_A[811]),
        .A_812(q_A[812]),
        .A_813(q_A[813]),
        .A_814(q_A[814]),
        .A_815(q_A[815]),
        .A_816(q_A[816]),
        .A_817(q_A[817]),
        .A_818(q_A[818]),
        .A_819(q_A[819]),
        .A_820(q_A[820]),
        .A_821(q_A[821]),
        .A_822(q_A[822]),
        .A_823(q_A[823]),
        .A_824(q_A[824]),
        .A_825(q_A[825]),
        .A_826(q_A[826]),
        .A_827(q_A[827]),
        .A_828(q_A[828]),
        .A_829(q_A[829]),
        .A_830(q_A[830]),
        .A_831(q_A[831]),
        .A_832(q_A[832]),
        .A_833(q_A[833]),
        .A_834(q_A[834]),
        .A_835(q_A[835]),
        .A_836(q_A[836]),
        .A_837(q_A[837]),
        .A_838(q_A[838]),
        .A_839(q_A[839]),
        .A_840(q_A[840]),
        .A_841(q_A[841]),
        .A_842(q_A[842]),
        .A_843(q_A[843]),
        .A_844(q_A[844]),
        .A_845(q_A[845]),
        .A_846(q_A[846]),
        .A_847(q_A[847]),
        .A_848(q_A[848]),
        .A_849(q_A[849]),
        .A_850(q_A[850]),
        .A_851(q_A[851]),
        .A_852(q_A[852]),
        .A_853(q_A[853]),
        .A_854(q_A[854]),
        .A_855(q_A[855]),
        .A_856(q_A[856]),
        .A_857(q_A[857]),
        .A_858(q_A[858]),
        .A_859(q_A[859]),
        .A_860(q_A[860]),
        .A_861(q_A[861]),
        .A_862(q_A[862]),
        .A_863(q_A[863]),
        .A_864(q_A[864]),
        .A_865(q_A[865]),
        .A_866(q_A[866]),
        .A_867(q_A[867]),
        .A_868(q_A[868]),
        .A_869(q_A[869]),
        .A_870(q_A[870]),
        .A_871(q_A[871]),
        .A_872(q_A[872]),
        .A_873(q_A[873]),
        .A_874(q_A[874]),
        .A_875(q_A[875]),
        .A_876(q_A[876]),
        .A_877(q_A[877]),
        .A_878(q_A[878]),
        .A_879(q_A[879]),
        .A_880(q_A[880]),
        .A_881(q_A[881]),
        .A_882(q_A[882]),
        .A_883(q_A[883]),
        .A_884(q_A[884]),
        .A_885(q_A[885]),
        .A_886(q_A[886]),
        .A_887(q_A[887]),
        .A_888(q_A[888]),
        .A_889(q_A[889]),
        .A_890(q_A[890]),
        .A_891(q_A[891]),
        .A_892(q_A[892]),
        .A_893(q_A[893]),
        .A_894(q_A[894]),
        .A_895(q_A[895]),
        .A_896(q_A[896]),
        .A_897(q_A[897]),
        .A_898(q_A[898]),
        .A_899(q_A[899]),
        .A_900(q_A[900]),
        .A_901(q_A[901]),
        .A_902(q_A[902]),
        .A_903(q_A[903]),
        .A_904(q_A[904]),
        .A_905(q_A[905]),
        .A_906(q_A[906]),
        .A_907(q_A[907]),
        .A_908(q_A[908]),
        .A_909(q_A[909]),
        .A_910(q_A[910]),
        .A_911(q_A[911]),
        .A_912(q_A[912]),
        .A_913(q_A[913]),
        .A_914(q_A[914]),
        .A_915(q_A[915]),
        .A_916(q_A[916]),
        .A_917(q_A[917]),
        .A_918(q_A[918]),
        .A_919(q_A[919]),
        .A_920(q_A[920]),
        .A_921(q_A[921]),
        .A_922(q_A[922]),
        .A_923(q_A[923]),
        .A_924(q_A[924]),
        .A_925(q_A[925]),
        .A_926(q_A[926]),
        .A_927(q_A[927]),
        .A_928(q_A[928]),
        .A_929(q_A[929]),
        .A_930(q_A[930]),
        .A_931(q_A[931]),
        .A_932(q_A[932]),
        .A_933(q_A[933]),
        .A_934(q_A[934]),
        .A_935(q_A[935]),
        .A_936(q_A[936]),
        .A_937(q_A[937]),
        .A_938(q_A[938]),
        .A_939(q_A[939]),
        .A_940(q_A[940]),
        .A_941(q_A[941]),
        .A_942(q_A[942]),
        .A_943(q_A[943]),
        .A_944(q_A[944]),
        .A_945(q_A[945]),
        .A_946(q_A[946]),
        .A_947(q_A[947]),
        .A_948(q_A[948]),
        .A_949(q_A[949]),
        .A_950(q_A[950]),
        .A_951(q_A[951]),
        .A_952(q_A[952]),
        .A_953(q_A[953]),
        .A_954(q_A[954]),
        .A_955(q_A[955]),
        .A_956(q_A[956]),
        .A_957(q_A[957]),
        .A_958(q_A[958]),
        .A_959(q_A[959]),
        .A_960(q_A[960]),
        .A_961(q_A[961]),
        .A_962(q_A[962]),
        .A_963(q_A[963]),
        .A_964(q_A[964]),
        .A_965(q_A[965]),
        .A_966(q_A[966]),
        .A_967(q_A[967]),
        .A_968(q_A[968]),
        .A_969(q_A[969]),
        .A_970(q_A[970]),
        .A_971(q_A[971]),
        .A_972(q_A[972]),
        .A_973(q_A[973]),
        .A_974(q_A[974]),
        .A_975(q_A[975]),
        .A_976(q_A[976]),
        .A_977(q_A[977]),
        .A_978(q_A[978]),
        .A_979(q_A[979]),
        .A_980(q_A[980]),
        .A_981(q_A[981]),
        .A_982(q_A[982]),
        .A_983(q_A[983]),
        .A_984(q_A[984]),
        .A_985(q_A[985]),
        .A_986(q_A[986]),
        .A_987(q_A[987]),
        .A_988(q_A[988]),
        .A_989(q_A[989]),
        .A_990(q_A[990]),
        .A_991(q_A[991]),
        .A_992(q_A[992]),
        .A_993(q_A[993]),
        .A_994(q_A[994]),
        .A_995(q_A[995]),
        .A_996(q_A[996]),
        .A_997(q_A[997]),
        .A_998(q_A[998]),
        .A_999(q_A[999]),
        .A_1000(q_A[1000]),
        .A_1001(q_A[1001]),
        .A_1002(q_A[1002]),
        .A_1003(q_A[1003]),
        .A_1004(q_A[1004]),
        .A_1005(q_A[1005]),
        .A_1006(q_A[1006]),
        .A_1007(q_A[1007]),
        .A_1008(q_A[1008]),
        .A_1009(q_A[1009]),
        .A_1010(q_A[1010]),
        .A_1011(q_A[1011]),
        .A_1012(q_A[1012]),
        .A_1013(q_A[1013]),
        .A_1014(q_A[1014]),
        .A_1015(q_A[1015]),
        .A_1016(q_A[1016]),
        .A_1017(q_A[1017]),
        .A_1018(q_A[1018]),
        .A_1019(q_A[1019]),
        .A_1020(q_A[1020]),
        .A_1021(q_A[1021]),
        .A_1022(q_A[1022]),
        .A_1023(q_A[1023]),
        .B_0(q_B[0]),
        .B_1(q_B[1]),
        .B_2(q_B[2]),
        .B_3(q_B[3]),
        .B_4(q_B[4]),
        .B_5(q_B[5]),
        .B_6(q_B[6]),
        .B_7(q_B[7]),
        .B_8(q_B[8]),
        .B_9(q_B[9]),
        .B_10(q_B[10]),
        .B_11(q_B[11]),
        .B_12(q_B[12]),
        .B_13(q_B[13]),
        .B_14(q_B[14]),
        .B_15(q_B[15]),
        .B_16(q_B[16]),
        .B_17(q_B[17]),
        .B_18(q_B[18]),
        .B_19(q_B[19]),
        .B_20(q_B[20]),
        .B_21(q_B[21]),
        .B_22(q_B[22]),
        .B_23(q_B[23]),
        .B_24(q_B[24]),
        .B_25(q_B[25]),
        .B_26(q_B[26]),
        .B_27(q_B[27]),
        .B_28(q_B[28]),
        .B_29(q_B[29]),
        .B_30(q_B[30]),
        .B_31(q_B[31]),
        .B_32(q_B[32]),
        .B_33(q_B[33]),
        .B_34(q_B[34]),
        .B_35(q_B[35]),
        .B_36(q_B[36]),
        .B_37(q_B[37]),
        .B_38(q_B[38]),
        .B_39(q_B[39]),
        .B_40(q_B[40]),
        .B_41(q_B[41]),
        .B_42(q_B[42]),
        .B_43(q_B[43]),
        .B_44(q_B[44]),
        .B_45(q_B[45]),
        .B_46(q_B[46]),
        .B_47(q_B[47]),
        .B_48(q_B[48]),
        .B_49(q_B[49]),
        .B_50(q_B[50]),
        .B_51(q_B[51]),
        .B_52(q_B[52]),
        .B_53(q_B[53]),
        .B_54(q_B[54]),
        .B_55(q_B[55]),
        .B_56(q_B[56]),
        .B_57(q_B[57]),
        .B_58(q_B[58]),
        .B_59(q_B[59]),
        .B_60(q_B[60]),
        .B_61(q_B[61]),
        .B_62(q_B[62]),
        .B_63(q_B[63]),
        .B_64(q_B[64]),
        .B_65(q_B[65]),
        .B_66(q_B[66]),
        .B_67(q_B[67]),
        .B_68(q_B[68]),
        .B_69(q_B[69]),
        .B_70(q_B[70]),
        .B_71(q_B[71]),
        .B_72(q_B[72]),
        .B_73(q_B[73]),
        .B_74(q_B[74]),
        .B_75(q_B[75]),
        .B_76(q_B[76]),
        .B_77(q_B[77]),
        .B_78(q_B[78]),
        .B_79(q_B[79]),
        .B_80(q_B[80]),
        .B_81(q_B[81]),
        .B_82(q_B[82]),
        .B_83(q_B[83]),
        .B_84(q_B[84]),
        .B_85(q_B[85]),
        .B_86(q_B[86]),
        .B_87(q_B[87]),
        .B_88(q_B[88]),
        .B_89(q_B[89]),
        .B_90(q_B[90]),
        .B_91(q_B[91]),
        .B_92(q_B[92]),
        .B_93(q_B[93]),
        .B_94(q_B[94]),
        .B_95(q_B[95]),
        .B_96(q_B[96]),
        .B_97(q_B[97]),
        .B_98(q_B[98]),
        .B_99(q_B[99]),
        .B_100(q_B[100]),
        .B_101(q_B[101]),
        .B_102(q_B[102]),
        .B_103(q_B[103]),
        .B_104(q_B[104]),
        .B_105(q_B[105]),
        .B_106(q_B[106]),
        .B_107(q_B[107]),
        .B_108(q_B[108]),
        .B_109(q_B[109]),
        .B_110(q_B[110]),
        .B_111(q_B[111]),
        .B_112(q_B[112]),
        .B_113(q_B[113]),
        .B_114(q_B[114]),
        .B_115(q_B[115]),
        .B_116(q_B[116]),
        .B_117(q_B[117]),
        .B_118(q_B[118]),
        .B_119(q_B[119]),
        .B_120(q_B[120]),
        .B_121(q_B[121]),
        .B_122(q_B[122]),
        .B_123(q_B[123]),
        .B_124(q_B[124]),
        .B_125(q_B[125]),
        .B_126(q_B[126]),
        .B_127(q_B[127]),
        .B_128(q_B[128]),
        .B_129(q_B[129]),
        .B_130(q_B[130]),
        .B_131(q_B[131]),
        .B_132(q_B[132]),
        .B_133(q_B[133]),
        .B_134(q_B[134]),
        .B_135(q_B[135]),
        .B_136(q_B[136]),
        .B_137(q_B[137]),
        .B_138(q_B[138]),
        .B_139(q_B[139]),
        .B_140(q_B[140]),
        .B_141(q_B[141]),
        .B_142(q_B[142]),
        .B_143(q_B[143]),
        .B_144(q_B[144]),
        .B_145(q_B[145]),
        .B_146(q_B[146]),
        .B_147(q_B[147]),
        .B_148(q_B[148]),
        .B_149(q_B[149]),
        .B_150(q_B[150]),
        .B_151(q_B[151]),
        .B_152(q_B[152]),
        .B_153(q_B[153]),
        .B_154(q_B[154]),
        .B_155(q_B[155]),
        .B_156(q_B[156]),
        .B_157(q_B[157]),
        .B_158(q_B[158]),
        .B_159(q_B[159]),
        .B_160(q_B[160]),
        .B_161(q_B[161]),
        .B_162(q_B[162]),
        .B_163(q_B[163]),
        .B_164(q_B[164]),
        .B_165(q_B[165]),
        .B_166(q_B[166]),
        .B_167(q_B[167]),
        .B_168(q_B[168]),
        .B_169(q_B[169]),
        .B_170(q_B[170]),
        .B_171(q_B[171]),
        .B_172(q_B[172]),
        .B_173(q_B[173]),
        .B_174(q_B[174]),
        .B_175(q_B[175]),
        .B_176(q_B[176]),
        .B_177(q_B[177]),
        .B_178(q_B[178]),
        .B_179(q_B[179]),
        .B_180(q_B[180]),
        .B_181(q_B[181]),
        .B_182(q_B[182]),
        .B_183(q_B[183]),
        .B_184(q_B[184]),
        .B_185(q_B[185]),
        .B_186(q_B[186]),
        .B_187(q_B[187]),
        .B_188(q_B[188]),
        .B_189(q_B[189]),
        .B_190(q_B[190]),
        .B_191(q_B[191]),
        .B_192(q_B[192]),
        .B_193(q_B[193]),
        .B_194(q_B[194]),
        .B_195(q_B[195]),
        .B_196(q_B[196]),
        .B_197(q_B[197]),
        .B_198(q_B[198]),
        .B_199(q_B[199]),
        .B_200(q_B[200]),
        .B_201(q_B[201]),
        .B_202(q_B[202]),
        .B_203(q_B[203]),
        .B_204(q_B[204]),
        .B_205(q_B[205]),
        .B_206(q_B[206]),
        .B_207(q_B[207]),
        .B_208(q_B[208]),
        .B_209(q_B[209]),
        .B_210(q_B[210]),
        .B_211(q_B[211]),
        .B_212(q_B[212]),
        .B_213(q_B[213]),
        .B_214(q_B[214]),
        .B_215(q_B[215]),
        .B_216(q_B[216]),
        .B_217(q_B[217]),
        .B_218(q_B[218]),
        .B_219(q_B[219]),
        .B_220(q_B[220]),
        .B_221(q_B[221]),
        .B_222(q_B[222]),
        .B_223(q_B[223]),
        .B_224(q_B[224]),
        .B_225(q_B[225]),
        .B_226(q_B[226]),
        .B_227(q_B[227]),
        .B_228(q_B[228]),
        .B_229(q_B[229]),
        .B_230(q_B[230]),
        .B_231(q_B[231]),
        .B_232(q_B[232]),
        .B_233(q_B[233]),
        .B_234(q_B[234]),
        .B_235(q_B[235]),
        .B_236(q_B[236]),
        .B_237(q_B[237]),
        .B_238(q_B[238]),
        .B_239(q_B[239]),
        .B_240(q_B[240]),
        .B_241(q_B[241]),
        .B_242(q_B[242]),
        .B_243(q_B[243]),
        .B_244(q_B[244]),
        .B_245(q_B[245]),
        .B_246(q_B[246]),
        .B_247(q_B[247]),
        .B_248(q_B[248]),
        .B_249(q_B[249]),
        .B_250(q_B[250]),
        .B_251(q_B[251]),
        .B_252(q_B[252]),
        .B_253(q_B[253]),
        .B_254(q_B[254]),
        .B_255(q_B[255]),
        .B_256(q_B[256]),
        .B_257(q_B[257]),
        .B_258(q_B[258]),
        .B_259(q_B[259]),
        .B_260(q_B[260]),
        .B_261(q_B[261]),
        .B_262(q_B[262]),
        .B_263(q_B[263]),
        .B_264(q_B[264]),
        .B_265(q_B[265]),
        .B_266(q_B[266]),
        .B_267(q_B[267]),
        .B_268(q_B[268]),
        .B_269(q_B[269]),
        .B_270(q_B[270]),
        .B_271(q_B[271]),
        .B_272(q_B[272]),
        .B_273(q_B[273]),
        .B_274(q_B[274]),
        .B_275(q_B[275]),
        .B_276(q_B[276]),
        .B_277(q_B[277]),
        .B_278(q_B[278]),
        .B_279(q_B[279]),
        .B_280(q_B[280]),
        .B_281(q_B[281]),
        .B_282(q_B[282]),
        .B_283(q_B[283]),
        .B_284(q_B[284]),
        .B_285(q_B[285]),
        .B_286(q_B[286]),
        .B_287(q_B[287]),
        .B_288(q_B[288]),
        .B_289(q_B[289]),
        .B_290(q_B[290]),
        .B_291(q_B[291]),
        .B_292(q_B[292]),
        .B_293(q_B[293]),
        .B_294(q_B[294]),
        .B_295(q_B[295]),
        .B_296(q_B[296]),
        .B_297(q_B[297]),
        .B_298(q_B[298]),
        .B_299(q_B[299]),
        .B_300(q_B[300]),
        .B_301(q_B[301]),
        .B_302(q_B[302]),
        .B_303(q_B[303]),
        .B_304(q_B[304]),
        .B_305(q_B[305]),
        .B_306(q_B[306]),
        .B_307(q_B[307]),
        .B_308(q_B[308]),
        .B_309(q_B[309]),
        .B_310(q_B[310]),
        .B_311(q_B[311]),
        .B_312(q_B[312]),
        .B_313(q_B[313]),
        .B_314(q_B[314]),
        .B_315(q_B[315]),
        .B_316(q_B[316]),
        .B_317(q_B[317]),
        .B_318(q_B[318]),
        .B_319(q_B[319]),
        .B_320(q_B[320]),
        .B_321(q_B[321]),
        .B_322(q_B[322]),
        .B_323(q_B[323]),
        .B_324(q_B[324]),
        .B_325(q_B[325]),
        .B_326(q_B[326]),
        .B_327(q_B[327]),
        .B_328(q_B[328]),
        .B_329(q_B[329]),
        .B_330(q_B[330]),
        .B_331(q_B[331]),
        .B_332(q_B[332]),
        .B_333(q_B[333]),
        .B_334(q_B[334]),
        .B_335(q_B[335]),
        .B_336(q_B[336]),
        .B_337(q_B[337]),
        .B_338(q_B[338]),
        .B_339(q_B[339]),
        .B_340(q_B[340]),
        .B_341(q_B[341]),
        .B_342(q_B[342]),
        .B_343(q_B[343]),
        .B_344(q_B[344]),
        .B_345(q_B[345]),
        .B_346(q_B[346]),
        .B_347(q_B[347]),
        .B_348(q_B[348]),
        .B_349(q_B[349]),
        .B_350(q_B[350]),
        .B_351(q_B[351]),
        .B_352(q_B[352]),
        .B_353(q_B[353]),
        .B_354(q_B[354]),
        .B_355(q_B[355]),
        .B_356(q_B[356]),
        .B_357(q_B[357]),
        .B_358(q_B[358]),
        .B_359(q_B[359]),
        .B_360(q_B[360]),
        .B_361(q_B[361]),
        .B_362(q_B[362]),
        .B_363(q_B[363]),
        .B_364(q_B[364]),
        .B_365(q_B[365]),
        .B_366(q_B[366]),
        .B_367(q_B[367]),
        .B_368(q_B[368]),
        .B_369(q_B[369]),
        .B_370(q_B[370]),
        .B_371(q_B[371]),
        .B_372(q_B[372]),
        .B_373(q_B[373]),
        .B_374(q_B[374]),
        .B_375(q_B[375]),
        .B_376(q_B[376]),
        .B_377(q_B[377]),
        .B_378(q_B[378]),
        .B_379(q_B[379]),
        .B_380(q_B[380]),
        .B_381(q_B[381]),
        .B_382(q_B[382]),
        .B_383(q_B[383]),
        .B_384(q_B[384]),
        .B_385(q_B[385]),
        .B_386(q_B[386]),
        .B_387(q_B[387]),
        .B_388(q_B[388]),
        .B_389(q_B[389]),
        .B_390(q_B[390]),
        .B_391(q_B[391]),
        .B_392(q_B[392]),
        .B_393(q_B[393]),
        .B_394(q_B[394]),
        .B_395(q_B[395]),
        .B_396(q_B[396]),
        .B_397(q_B[397]),
        .B_398(q_B[398]),
        .B_399(q_B[399]),
        .B_400(q_B[400]),
        .B_401(q_B[401]),
        .B_402(q_B[402]),
        .B_403(q_B[403]),
        .B_404(q_B[404]),
        .B_405(q_B[405]),
        .B_406(q_B[406]),
        .B_407(q_B[407]),
        .B_408(q_B[408]),
        .B_409(q_B[409]),
        .B_410(q_B[410]),
        .B_411(q_B[411]),
        .B_412(q_B[412]),
        .B_413(q_B[413]),
        .B_414(q_B[414]),
        .B_415(q_B[415]),
        .B_416(q_B[416]),
        .B_417(q_B[417]),
        .B_418(q_B[418]),
        .B_419(q_B[419]),
        .B_420(q_B[420]),
        .B_421(q_B[421]),
        .B_422(q_B[422]),
        .B_423(q_B[423]),
        .B_424(q_B[424]),
        .B_425(q_B[425]),
        .B_426(q_B[426]),
        .B_427(q_B[427]),
        .B_428(q_B[428]),
        .B_429(q_B[429]),
        .B_430(q_B[430]),
        .B_431(q_B[431]),
        .B_432(q_B[432]),
        .B_433(q_B[433]),
        .B_434(q_B[434]),
        .B_435(q_B[435]),
        .B_436(q_B[436]),
        .B_437(q_B[437]),
        .B_438(q_B[438]),
        .B_439(q_B[439]),
        .B_440(q_B[440]),
        .B_441(q_B[441]),
        .B_442(q_B[442]),
        .B_443(q_B[443]),
        .B_444(q_B[444]),
        .B_445(q_B[445]),
        .B_446(q_B[446]),
        .B_447(q_B[447]),
        .B_448(q_B[448]),
        .B_449(q_B[449]),
        .B_450(q_B[450]),
        .B_451(q_B[451]),
        .B_452(q_B[452]),
        .B_453(q_B[453]),
        .B_454(q_B[454]),
        .B_455(q_B[455]),
        .B_456(q_B[456]),
        .B_457(q_B[457]),
        .B_458(q_B[458]),
        .B_459(q_B[459]),
        .B_460(q_B[460]),
        .B_461(q_B[461]),
        .B_462(q_B[462]),
        .B_463(q_B[463]),
        .B_464(q_B[464]),
        .B_465(q_B[465]),
        .B_466(q_B[466]),
        .B_467(q_B[467]),
        .B_468(q_B[468]),
        .B_469(q_B[469]),
        .B_470(q_B[470]),
        .B_471(q_B[471]),
        .B_472(q_B[472]),
        .B_473(q_B[473]),
        .B_474(q_B[474]),
        .B_475(q_B[475]),
        .B_476(q_B[476]),
        .B_477(q_B[477]),
        .B_478(q_B[478]),
        .B_479(q_B[479]),
        .B_480(q_B[480]),
        .B_481(q_B[481]),
        .B_482(q_B[482]),
        .B_483(q_B[483]),
        .B_484(q_B[484]),
        .B_485(q_B[485]),
        .B_486(q_B[486]),
        .B_487(q_B[487]),
        .B_488(q_B[488]),
        .B_489(q_B[489]),
        .B_490(q_B[490]),
        .B_491(q_B[491]),
        .B_492(q_B[492]),
        .B_493(q_B[493]),
        .B_494(q_B[494]),
        .B_495(q_B[495]),
        .B_496(q_B[496]),
        .B_497(q_B[497]),
        .B_498(q_B[498]),
        .B_499(q_B[499]),
        .B_500(q_B[500]),
        .B_501(q_B[501]),
        .B_502(q_B[502]),
        .B_503(q_B[503]),
        .B_504(q_B[504]),
        .B_505(q_B[505]),
        .B_506(q_B[506]),
        .B_507(q_B[507]),
        .B_508(q_B[508]),
        .B_509(q_B[509]),
        .B_510(q_B[510]),
        .B_511(q_B[511]),
        .B_512(q_B[512]),
        .B_513(q_B[513]),
        .B_514(q_B[514]),
        .B_515(q_B[515]),
        .B_516(q_B[516]),
        .B_517(q_B[517]),
        .B_518(q_B[518]),
        .B_519(q_B[519]),
        .B_520(q_B[520]),
        .B_521(q_B[521]),
        .B_522(q_B[522]),
        .B_523(q_B[523]),
        .B_524(q_B[524]),
        .B_525(q_B[525]),
        .B_526(q_B[526]),
        .B_527(q_B[527]),
        .B_528(q_B[528]),
        .B_529(q_B[529]),
        .B_530(q_B[530]),
        .B_531(q_B[531]),
        .B_532(q_B[532]),
        .B_533(q_B[533]),
        .B_534(q_B[534]),
        .B_535(q_B[535]),
        .B_536(q_B[536]),
        .B_537(q_B[537]),
        .B_538(q_B[538]),
        .B_539(q_B[539]),
        .B_540(q_B[540]),
        .B_541(q_B[541]),
        .B_542(q_B[542]),
        .B_543(q_B[543]),
        .B_544(q_B[544]),
        .B_545(q_B[545]),
        .B_546(q_B[546]),
        .B_547(q_B[547]),
        .B_548(q_B[548]),
        .B_549(q_B[549]),
        .B_550(q_B[550]),
        .B_551(q_B[551]),
        .B_552(q_B[552]),
        .B_553(q_B[553]),
        .B_554(q_B[554]),
        .B_555(q_B[555]),
        .B_556(q_B[556]),
        .B_557(q_B[557]),
        .B_558(q_B[558]),
        .B_559(q_B[559]),
        .B_560(q_B[560]),
        .B_561(q_B[561]),
        .B_562(q_B[562]),
        .B_563(q_B[563]),
        .B_564(q_B[564]),
        .B_565(q_B[565]),
        .B_566(q_B[566]),
        .B_567(q_B[567]),
        .B_568(q_B[568]),
        .B_569(q_B[569]),
        .B_570(q_B[570]),
        .B_571(q_B[571]),
        .B_572(q_B[572]),
        .B_573(q_B[573]),
        .B_574(q_B[574]),
        .B_575(q_B[575]),
        .B_576(q_B[576]),
        .B_577(q_B[577]),
        .B_578(q_B[578]),
        .B_579(q_B[579]),
        .B_580(q_B[580]),
        .B_581(q_B[581]),
        .B_582(q_B[582]),
        .B_583(q_B[583]),
        .B_584(q_B[584]),
        .B_585(q_B[585]),
        .B_586(q_B[586]),
        .B_587(q_B[587]),
        .B_588(q_B[588]),
        .B_589(q_B[589]),
        .B_590(q_B[590]),
        .B_591(q_B[591]),
        .B_592(q_B[592]),
        .B_593(q_B[593]),
        .B_594(q_B[594]),
        .B_595(q_B[595]),
        .B_596(q_B[596]),
        .B_597(q_B[597]),
        .B_598(q_B[598]),
        .B_599(q_B[599]),
        .B_600(q_B[600]),
        .B_601(q_B[601]),
        .B_602(q_B[602]),
        .B_603(q_B[603]),
        .B_604(q_B[604]),
        .B_605(q_B[605]),
        .B_606(q_B[606]),
        .B_607(q_B[607]),
        .B_608(q_B[608]),
        .B_609(q_B[609]),
        .B_610(q_B[610]),
        .B_611(q_B[611]),
        .B_612(q_B[612]),
        .B_613(q_B[613]),
        .B_614(q_B[614]),
        .B_615(q_B[615]),
        .B_616(q_B[616]),
        .B_617(q_B[617]),
        .B_618(q_B[618]),
        .B_619(q_B[619]),
        .B_620(q_B[620]),
        .B_621(q_B[621]),
        .B_622(q_B[622]),
        .B_623(q_B[623]),
        .B_624(q_B[624]),
        .B_625(q_B[625]),
        .B_626(q_B[626]),
        .B_627(q_B[627]),
        .B_628(q_B[628]),
        .B_629(q_B[629]),
        .B_630(q_B[630]),
        .B_631(q_B[631]),
        .B_632(q_B[632]),
        .B_633(q_B[633]),
        .B_634(q_B[634]),
        .B_635(q_B[635]),
        .B_636(q_B[636]),
        .B_637(q_B[637]),
        .B_638(q_B[638]),
        .B_639(q_B[639]),
        .B_640(q_B[640]),
        .B_641(q_B[641]),
        .B_642(q_B[642]),
        .B_643(q_B[643]),
        .B_644(q_B[644]),
        .B_645(q_B[645]),
        .B_646(q_B[646]),
        .B_647(q_B[647]),
        .B_648(q_B[648]),
        .B_649(q_B[649]),
        .B_650(q_B[650]),
        .B_651(q_B[651]),
        .B_652(q_B[652]),
        .B_653(q_B[653]),
        .B_654(q_B[654]),
        .B_655(q_B[655]),
        .B_656(q_B[656]),
        .B_657(q_B[657]),
        .B_658(q_B[658]),
        .B_659(q_B[659]),
        .B_660(q_B[660]),
        .B_661(q_B[661]),
        .B_662(q_B[662]),
        .B_663(q_B[663]),
        .B_664(q_B[664]),
        .B_665(q_B[665]),
        .B_666(q_B[666]),
        .B_667(q_B[667]),
        .B_668(q_B[668]),
        .B_669(q_B[669]),
        .B_670(q_B[670]),
        .B_671(q_B[671]),
        .B_672(q_B[672]),
        .B_673(q_B[673]),
        .B_674(q_B[674]),
        .B_675(q_B[675]),
        .B_676(q_B[676]),
        .B_677(q_B[677]),
        .B_678(q_B[678]),
        .B_679(q_B[679]),
        .B_680(q_B[680]),
        .B_681(q_B[681]),
        .B_682(q_B[682]),
        .B_683(q_B[683]),
        .B_684(q_B[684]),
        .B_685(q_B[685]),
        .B_686(q_B[686]),
        .B_687(q_B[687]),
        .B_688(q_B[688]),
        .B_689(q_B[689]),
        .B_690(q_B[690]),
        .B_691(q_B[691]),
        .B_692(q_B[692]),
        .B_693(q_B[693]),
        .B_694(q_B[694]),
        .B_695(q_B[695]),
        .B_696(q_B[696]),
        .B_697(q_B[697]),
        .B_698(q_B[698]),
        .B_699(q_B[699]),
        .B_700(q_B[700]),
        .B_701(q_B[701]),
        .B_702(q_B[702]),
        .B_703(q_B[703]),
        .B_704(q_B[704]),
        .B_705(q_B[705]),
        .B_706(q_B[706]),
        .B_707(q_B[707]),
        .B_708(q_B[708]),
        .B_709(q_B[709]),
        .B_710(q_B[710]),
        .B_711(q_B[711]),
        .B_712(q_B[712]),
        .B_713(q_B[713]),
        .B_714(q_B[714]),
        .B_715(q_B[715]),
        .B_716(q_B[716]),
        .B_717(q_B[717]),
        .B_718(q_B[718]),
        .B_719(q_B[719]),
        .B_720(q_B[720]),
        .B_721(q_B[721]),
        .B_722(q_B[722]),
        .B_723(q_B[723]),
        .B_724(q_B[724]),
        .B_725(q_B[725]),
        .B_726(q_B[726]),
        .B_727(q_B[727]),
        .B_728(q_B[728]),
        .B_729(q_B[729]),
        .B_730(q_B[730]),
        .B_731(q_B[731]),
        .B_732(q_B[732]),
        .B_733(q_B[733]),
        .B_734(q_B[734]),
        .B_735(q_B[735]),
        .B_736(q_B[736]),
        .B_737(q_B[737]),
        .B_738(q_B[738]),
        .B_739(q_B[739]),
        .B_740(q_B[740]),
        .B_741(q_B[741]),
        .B_742(q_B[742]),
        .B_743(q_B[743]),
        .B_744(q_B[744]),
        .B_745(q_B[745]),
        .B_746(q_B[746]),
        .B_747(q_B[747]),
        .B_748(q_B[748]),
        .B_749(q_B[749]),
        .B_750(q_B[750]),
        .B_751(q_B[751]),
        .B_752(q_B[752]),
        .B_753(q_B[753]),
        .B_754(q_B[754]),
        .B_755(q_B[755]),
        .B_756(q_B[756]),
        .B_757(q_B[757]),
        .B_758(q_B[758]),
        .B_759(q_B[759]),
        .B_760(q_B[760]),
        .B_761(q_B[761]),
        .B_762(q_B[762]),
        .B_763(q_B[763]),
        .B_764(q_B[764]),
        .B_765(q_B[765]),
        .B_766(q_B[766]),
        .B_767(q_B[767]),
        .B_768(q_B[768]),
        .B_769(q_B[769]),
        .B_770(q_B[770]),
        .B_771(q_B[771]),
        .B_772(q_B[772]),
        .B_773(q_B[773]),
        .B_774(q_B[774]),
        .B_775(q_B[775]),
        .B_776(q_B[776]),
        .B_777(q_B[777]),
        .B_778(q_B[778]),
        .B_779(q_B[779]),
        .B_780(q_B[780]),
        .B_781(q_B[781]),
        .B_782(q_B[782]),
        .B_783(q_B[783]),
        .B_784(q_B[784]),
        .B_785(q_B[785]),
        .B_786(q_B[786]),
        .B_787(q_B[787]),
        .B_788(q_B[788]),
        .B_789(q_B[789]),
        .B_790(q_B[790]),
        .B_791(q_B[791]),
        .B_792(q_B[792]),
        .B_793(q_B[793]),
        .B_794(q_B[794]),
        .B_795(q_B[795]),
        .B_796(q_B[796]),
        .B_797(q_B[797]),
        .B_798(q_B[798]),
        .B_799(q_B[799]),
        .B_800(q_B[800]),
        .B_801(q_B[801]),
        .B_802(q_B[802]),
        .B_803(q_B[803]),
        .B_804(q_B[804]),
        .B_805(q_B[805]),
        .B_806(q_B[806]),
        .B_807(q_B[807]),
        .B_808(q_B[808]),
        .B_809(q_B[809]),
        .B_810(q_B[810]),
        .B_811(q_B[811]),
        .B_812(q_B[812]),
        .B_813(q_B[813]),
        .B_814(q_B[814]),
        .B_815(q_B[815]),
        .B_816(q_B[816]),
        .B_817(q_B[817]),
        .B_818(q_B[818]),
        .B_819(q_B[819]),
        .B_820(q_B[820]),
        .B_821(q_B[821]),
        .B_822(q_B[822]),
        .B_823(q_B[823]),
        .B_824(q_B[824]),
        .B_825(q_B[825]),
        .B_826(q_B[826]),
        .B_827(q_B[827]),
        .B_828(q_B[828]),
        .B_829(q_B[829]),
        .B_830(q_B[830]),
        .B_831(q_B[831]),
        .B_832(q_B[832]),
        .B_833(q_B[833]),
        .B_834(q_B[834]),
        .B_835(q_B[835]),
        .B_836(q_B[836]),
        .B_837(q_B[837]),
        .B_838(q_B[838]),
        .B_839(q_B[839]),
        .B_840(q_B[840]),
        .B_841(q_B[841]),
        .B_842(q_B[842]),
        .B_843(q_B[843]),
        .B_844(q_B[844]),
        .B_845(q_B[845]),
        .B_846(q_B[846]),
        .B_847(q_B[847]),
        .B_848(q_B[848]),
        .B_849(q_B[849]),
        .B_850(q_B[850]),
        .B_851(q_B[851]),
        .B_852(q_B[852]),
        .B_853(q_B[853]),
        .B_854(q_B[854]),
        .B_855(q_B[855]),
        .B_856(q_B[856]),
        .B_857(q_B[857]),
        .B_858(q_B[858]),
        .B_859(q_B[859]),
        .B_860(q_B[860]),
        .B_861(q_B[861]),
        .B_862(q_B[862]),
        .B_863(q_B[863]),
        .B_864(q_B[864]),
        .B_865(q_B[865]),
        .B_866(q_B[866]),
        .B_867(q_B[867]),
        .B_868(q_B[868]),
        .B_869(q_B[869]),
        .B_870(q_B[870]),
        .B_871(q_B[871]),
        .B_872(q_B[872]),
        .B_873(q_B[873]),
        .B_874(q_B[874]),
        .B_875(q_B[875]),
        .B_876(q_B[876]),
        .B_877(q_B[877]),
        .B_878(q_B[878]),
        .B_879(q_B[879]),
        .B_880(q_B[880]),
        .B_881(q_B[881]),
        .B_882(q_B[882]),
        .B_883(q_B[883]),
        .B_884(q_B[884]),
        .B_885(q_B[885]),
        .B_886(q_B[886]),
        .B_887(q_B[887]),
        .B_888(q_B[888]),
        .B_889(q_B[889]),
        .B_890(q_B[890]),
        .B_891(q_B[891]),
        .B_892(q_B[892]),
        .B_893(q_B[893]),
        .B_894(q_B[894]),
        .B_895(q_B[895]),
        .B_896(q_B[896]),
        .B_897(q_B[897]),
        .B_898(q_B[898]),
        .B_899(q_B[899]),
        .B_900(q_B[900]),
        .B_901(q_B[901]),
        .B_902(q_B[902]),
        .B_903(q_B[903]),
        .B_904(q_B[904]),
        .B_905(q_B[905]),
        .B_906(q_B[906]),
        .B_907(q_B[907]),
        .B_908(q_B[908]),
        .B_909(q_B[909]),
        .B_910(q_B[910]),
        .B_911(q_B[911]),
        .B_912(q_B[912]),
        .B_913(q_B[913]),
        .B_914(q_B[914]),
        .B_915(q_B[915]),
        .B_916(q_B[916]),
        .B_917(q_B[917]),
        .B_918(q_B[918]),
        .B_919(q_B[919]),
        .B_920(q_B[920]),
        .B_921(q_B[921]),
        .B_922(q_B[922]),
        .B_923(q_B[923]),
        .B_924(q_B[924]),
        .B_925(q_B[925]),
        .B_926(q_B[926]),
        .B_927(q_B[927]),
        .B_928(q_B[928]),
        .B_929(q_B[929]),
        .B_930(q_B[930]),
        .B_931(q_B[931]),
        .B_932(q_B[932]),
        .B_933(q_B[933]),
        .B_934(q_B[934]),
        .B_935(q_B[935]),
        .B_936(q_B[936]),
        .B_937(q_B[937]),
        .B_938(q_B[938]),
        .B_939(q_B[939]),
        .B_940(q_B[940]),
        .B_941(q_B[941]),
        .B_942(q_B[942]),
        .B_943(q_B[943]),
        .B_944(q_B[944]),
        .B_945(q_B[945]),
        .B_946(q_B[946]),
        .B_947(q_B[947]),
        .B_948(q_B[948]),
        .B_949(q_B[949]),
        .B_950(q_B[950]),
        .B_951(q_B[951]),
        .B_952(q_B[952]),
        .B_953(q_B[953]),
        .B_954(q_B[954]),
        .B_955(q_B[955]),
        .B_956(q_B[956]),
        .B_957(q_B[957]),
        .B_958(q_B[958]),
        .B_959(q_B[959]),
        .B_960(q_B[960]),
        .B_961(q_B[961]),
        .B_962(q_B[962]),
        .B_963(q_B[963]),
        .B_964(q_B[964]),
        .B_965(q_B[965]),
        .B_966(q_B[966]),
        .B_967(q_B[967]),
        .B_968(q_B[968]),
        .B_969(q_B[969]),
        .B_970(q_B[970]),
        .B_971(q_B[971]),
        .B_972(q_B[972]),
        .B_973(q_B[973]),
        .B_974(q_B[974]),
        .B_975(q_B[975]),
        .B_976(q_B[976]),
        .B_977(q_B[977]),
        .B_978(q_B[978]),
        .B_979(q_B[979]),
        .B_980(q_B[980]),
        .B_981(q_B[981]),
        .B_982(q_B[982]),
        .B_983(q_B[983]),
        .B_984(q_B[984]),
        .B_985(q_B[985]),
        .B_986(q_B[986]),
        .B_987(q_B[987]),
        .B_988(q_B[988]),
        .B_989(q_B[989]),
        .B_990(q_B[990]),
        .B_991(q_B[991]),
        .B_992(q_B[992]),
        .B_993(q_B[993]),
        .B_994(q_B[994]),
        .B_995(q_B[995]),
        .B_996(q_B[996]),
        .B_997(q_B[997]),
        .B_998(q_B[998]),
        .B_999(q_B[999]),
        .B_1000(q_B[1000]),
        .B_1001(q_B[1001]),
        .B_1002(q_B[1002]),
        .B_1003(q_B[1003]),
        .B_1004(q_B[1004]),
        .B_1005(q_B[1005]),
        .B_1006(q_B[1006]),
        .B_1007(q_B[1007]),
        .B_1008(q_B[1008]),
        .B_1009(q_B[1009]),
        .B_1010(q_B[1010]),
        .B_1011(q_B[1011]),
        .B_1012(q_B[1012]),
        .B_1013(q_B[1013]),
        .B_1014(q_B[1014]),
        .B_1015(q_B[1015]),
        .B_1016(q_B[1016]),
        .B_1017(q_B[1017]),
        .B_1018(q_B[1018]),
        .B_1019(q_B[1019]),
        .B_1020(q_B[1020]),
        .B_1021(q_B[1021]),
        .B_1022(q_B[1022]),
        .B_1023(q_B[1023])
    );


    // OUTPUT CONTROL
    control_out out_ctrl_inst (
        .clk(clk_out1), .reset(reset), 
        .ap_done(ap_done),
        .hls_result(hls_result), .hls_opcode(hls_opcode),
        .tx_busy(tx_busy),
        .tx_start(core_tx_start), .tx_data(core_tx_data),
        .disp_data(disp_data), .disp_opcode(disp_opcode)
    );

    // UART & DISPLAY
    uart_basic #(.CLK_FREQUENCY_RX(100000000)) uart_inst (
        .clk_rx(clk_out1), .reset_rx(reset), .rx(rx), 
        .rx_data(rx_data), .rx_ready(rx_ready),
        .clk_tx(clk_out1), .reset_tx(reset), .tx(tx), 
        .tx_start(core_tx_start), .tx_data(core_tx_data), 
        .tx_busy(tx_busy)
    );

    display_interface disp_inst (
        .clk(clk_out1), .reset(reset), 
        .data_in(disp_data), .opcode(disp_opcode),
        .an(an), .seg(seg), .dp(dp)
    );
    /*
    ila_0 my_ila (
        .clk(clk_out1),
        .probe0(ap_start),
        .probe1(ap_done),
        .probe2(hls_opcode),
        .probe3(hls_result) 
    );
    */
endmodule